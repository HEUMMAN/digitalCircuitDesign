library verilog;
use verilog.vl_types.all;
entity structural_mux_vlg_check_tst is
    port(
        \out\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end structural_mux_vlg_check_tst;
