library verilog;
use verilog.vl_types.all;
entity structural_mux_vlg_vec_tst is
end structural_mux_vlg_vec_tst;
