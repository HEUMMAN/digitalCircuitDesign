library verilog;
use verilog.vl_types.all;
entity DUT_TEST_tb is
end DUT_TEST_tb;
